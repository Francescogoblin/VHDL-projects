sdvhbsdjknsdjc
