library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-- andiamo a spezzare il processo combinatorio più lungo, così che il tempo di propagazione totale è 15ns


