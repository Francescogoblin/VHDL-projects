library IEEE;
	use IEEE.STD_LOGIC_1164.ALL;

entity ff_d is
	Port(
		reset	: in  std_logic;
		clk		: in  std_logic;

		d 	        : in  std_logic;
		q 	        : out std_logic
	);
end ff_d;

architecture Behavioral of ff_d is
	
	

begin

	
end Behavioral;
