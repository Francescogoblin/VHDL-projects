
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-- Latenza= 1 ciclo di clock = Tclk.  
-- Scelgo il tempo di clock minimo (che mi darà la frequenza massima) sapendo che non ha senso "riaprire il cancello" se la logica non ha ancora elaborato un risultato. Quindi Tclk=Tpd= 22ns
-- Throughput del sistema --> dipende dal tempo di clock. In questo caso sarà 1/Tclk = 45 Mhz 
-- Con un clock a 45MHz il throughput è 45MHz * 32bit al secondo = 45MHz * 4Byte al secondo = 1440 MBit/sec 

entity Esercizio2 is
  Port(
    input_a : in std_logic_vector ( 31 DOWNTO 0) ;
    input_b : in std_logic_vector ( 31 DOWNTO 0) ;
    input_c : in std_logic_vector ( 31 DOWNTO 0) ;
    clk     : in std_logic;
    reset	: in std_logic;
	  
    result  : out std_logic_vector ( 31 DOWNTO 0)
  );
end Esercizio2;
-----------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------
	
  Architecture Behavioral of Esercizio2 is 
  
    component multiplier is
	Port (
	input_a			: in unsigned(31 DOWNTO 0);
	input_b			: in unsigned(31 DOWNTO 0);
	result			: out unsigned(31 DOWNTO 0)
	);
    end component;
    
    component adder is
	Port (
	input_a			: in unsigned(31 DOWNTO 0);
	input_b			: in unsigned(31 DOWNTO 0);
	result			: out unsigned(31 DOWNTO 0)
	);
    end component;

    signal out_mul   : unsigned(31 DOWNTO 0);
	signal out_adder : unsigned(31 DOWNTO 0);

-----------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------

    begin

    MULTIPLIER_INST : multiplier
      Port map ( 
          input_a   => unsigned(input_a),
	      input_b	=> unsigned(input_b),
	      result	=> out_mul
      );
      
    ADDER_INST : adder
      Port map ( 
          input_a   => unsigned(input_c),
	      input_b	=> out_mul
	      result	=> out_adder -- out adder ora è ancora unsigned
      );

		-- fin qui tutto praticamente uguale a prima , cambia solo che ora ho un signal in più a cui collegare l'uscita dell'adder
		-- ora vado a fare il process per instanziare il registro
		process ( clk  , reset ) 
		begin
				if reset = '1' then
					result <= (Others => '0');
				end if;
					
				if rising_edge(clk) = '1' then
					result <= std_logic_vector(out_add);
				end if;
		end process;
      
 end Behavioral;   
    
