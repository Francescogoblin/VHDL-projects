library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ShiftRegisterSIPO is
	
Generic(
SR_WIDTH :integer:= 4
); 
Port(
reset    : in  std_logic;
clk      : in  std_logic;
data_in  : in  std_logic;
data_out : out std_logic_vector(SR_WIDTH-1 DOWNTO 0)
);     
end ShiftRegisterSIPO;


architecture Behavioral of ShiftRegisterSIPO is
	
	component ff_d is
    	Port(
			reset_ff	: in std_logic;
			clk_ff    : in std_logic;
			d 		: in std_logic;
			q 		: out std_logic
		);  
	end component;
	   
	signal n : std_logic_vector(3 DOWNTO 0);

begin
	if SR_WIDTH = 0 then
		
    	report "Errore: STD è uguale a 1" severity error;
	
	elsif SR_WIDTH > 0 then
	
	ff_d_inst_0 : ff_d                                                          --INSTANZA INIZIALE
    	Port Map (
        	reset_ff => reset,
            clk_ff   => clk,
        	d        => data_in,
       	    q        => n(0)
        );
            
   	LOOP_GEN  : for I in 0 to SR_WIDTH-2 generate                                 --INIZIO DEL LOOP
        
    ff_d_inst_i : ff_d
		Port Map (
        	reset_ff => reset,
            clk_ff   => clk,
        	d        => n(I),
        	q        => n(I+1)
        );
               
    end generate;
    	
	data_out <= n;

	end if;
                
end Behavioral;

