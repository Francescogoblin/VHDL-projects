--codice
